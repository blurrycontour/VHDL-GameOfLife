
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use ieee.std_logic_unsigned.all;


entity GoL is 
port
(	
	clr:in std_logic;
	hsync : out std_logic;
	vsync : out std_logic;
	clk_50 : in std_logic;
	red : out std_logic;
	green : out std_logic;
	blue : out std_logic;
	navy : out std_logic
	
	--hc : out std_logic_vector(9 downto 0);
	--vc : out std_logic_vector(9 downto 0);
	--btn : in std_logic_vector(3 downto 0);
	--vidon : out std_logic;
);
end GoL;



architecture GoL_a of GoL is

type Arr is array (23 downto 0, 31 downto 0) of integer;
type MArr is array (0 to 23, 0 to 31) of std_logic;
type arra is array (7 downto 0) of integer;
constant hpixels : std_logic_vector(9 downto 0) := "1100100000"; 
constant vlines : std_logic_vector(9 downto 0) := "1000001001";
constant hbp : std_logic_vector(9 downto 0) := "0010010000";
constant hfp : std_logic_vector(9 downto 0) := "1100010000";
constant vbp : std_logic_vector(9 downto 0) := "0000011111";
constant vfp : std_logic_vector(9 downto 0) := "0111111111";
signal clka : std_logic;
shared variable col,row :integer := 0;
shared variable decide : integer := 0;										  
--signal done : integer;
shared variable M : Arr :=((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
									(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

signal hcs,vcs : std_logic_vector(9 downto 0);
signal vsenable : std_logic;
signal clk : std_logic;
signal scalar : integer range 0 to 1;
signal scalara : integer range 0 to 25000000;
signal vidon ,done: std_logic;

--function neigh(K : integer;l : integer) return integer is
--variable counter: integer:= 0;
--begin
--	
--	if A(k-1)(l-1) = '1' then counter := counter + 1; end if;
--	if A(k-1)(l) = '1' then counter := counter + 1;end if;
--	if A(k-1)(l+1) = '1' then counter := counter + 1;end if;
--	if A(k)(l-1) = '1' then counter := counter + 1;end if;
--	if A(k)(l+1) = '1' then counter := counter + 1;end if;
--	if A(k+1)(l-1) = '1' then counter := counter + 1;end if;
--	if A(k+1)(l) = '1' then counter := counter + 1;end if;
--	if A(k+1)(l+1) = '1' then counter := counter + 1;end if;
--return counter;
--end function neigh;

--function state(bool1,bool2,bool3,bool4:boolean) return std_logic is
--variable ret : std_logic := '0';
--begin
--	if bool4 then 
--		ret := '1'; 
--	end if;
--	if bool3 then
--		ret := '1'; 
--	end if;
--	if bool1 then 
--		ret := '0'; 
--	end if;
--	if bool2 then 
--		ret := '0'; 
--	end if;
--
--return ret;
--end function state;


begin

	
	process( clk_50 , clr )
	begin
		if (clr = '0') then 
			clk <= '0';
			scalar <= 0;
		elsif(rising_edge(clk_50)) then 
			if (scalar < 1) then 
				scalar <= scalar + 1 ;
				clk <= '0';
			else
				scalar <= 0;
				clk <= '1';
			end if;
		end if;
	end process ;
	
	
	process( clk_50 , clr )
	begin
		if (clr = '0') then 
			clka <= '0';
			scalara <= 0;
		elsif(rising_edge(clk_50)) then 
			if (scalara < 25000000) then 
				scalara <= scalara + 1 ;
				clka <= '0';
			else
				scalara <= 0;
				clka <= '1';
			end if;
		end if;
	end process ;
	
	
	process(clk,clr,hcs)
	begin
		if clr = '0' then
			hcs <= "0000000000";
			col := to_integer(unsigned(hcs));
		elsif(clk'event and clk='1') then
			if hcs=hpixels-1 then 
				hcs <= "0000000000";
				col := to_integer(unsigned(hcs));
				vsenable <= '1';
			else
				hcs <= hcs + 1;
				col := to_integer(unsigned(hcs));
				vsenable <= '0';
			end if;
		end if;
	end process;	
			
	hsync <= '0' when hcs < 128 else '1';
	

	process(clk,clr,vcs)
	begin
		if clr = '0' then
			vcs <= "0000000000";
			row := to_integer(unsigned(vcs));
		elsif(clk'event and clk='1' and vsenable='1') then
			if vcs=vlines-1 then 
				vcs <= "0000000000";
				row := to_integer(unsigned(vcs));
			else
				vcs <= vcs + 1;
				row := to_integer(unsigned(vcs));
			end if;
		end if;
	end process;	
			
	vsync <= '0' when vcs < 2 else '1';
	
			
			
vidon <='1' when (((hcs < hfp) and (hcs >= hbp)) and 
						((vcs < vfp) and (vcs >= vbp)))  else '0';
						
	
	
--------------------------------------------------------------------------------------------	
	process(clka)
	
	variable n,cell : std_ulogic := '0';
	variable t : integer range 0 to 1 := 0 ;
	variable num: integer ;
	variable test : integer;
	variable boola,boolb,boolc,boold : boolean := false; 
	variable Ba,Bb,Bc,Bd : boolean := false;
	variable co : arra := (0,0,0,0,0,0,0,0);
	
	
	variable A : MArr :=(	('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','1','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','1','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','1','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','1','0','0','0','0','0','0','0','0','0','0','0'),
									('0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','0','1','0','0','0','0','0','0','0','0','0','0','0'),
									('0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','0','1','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','1','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','1','0','1','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','1','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','1','0','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0'),
									('0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','1','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','1','0','1','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
 
 variable B : MArr := (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
									('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
	begin
			
		if decide = 0 and rising_edge(clka) then 
		
			for I in 22 downto 1 loop 
				for J in 30 downto 1  loop				
					cell := A(I,J);				
							if (A(I-1,J-1) = '1') then 
								co(0) := 1; 
							else 
								co(0) := 0; 
							end if;
								if (A(I-1,J) = '1') then 
									co(1) := 1; 
								else 
									co(1) := 0;
								end if;
									if (A(I-1,J+1) = '1') then 
										co(2) := 1; 
									else 
										co(2) := 0;
									end if;
										if (A(I,J-1) = '1') then 
											co(3) := 1; 
										else 
											co(3) := 0;
										end if;
											if (A(I,J+1) = '1') then 
												co(4) := 1; 
											else 
												co(4) := 0;
											end if;
												if (A(I+1,J-1) = '1') then 
													co(5) := 1; 
												else 
													co(5) := 0;
												end if;
													if (A(I+1,J) = '1') then 
														co(6) := 1; 
													else 
														co(6) := 0;
													end if;
														if (A(I+1,J+1) = '1') then 
															co(7) := 1; 
														else 
															co(7) := 0;
														end if;				
																	M(I,J) := co(0)+co(1)+co(2)+co(3)+co(4)+co(5)+co(6)+co(7);
																		boola := ((M(I,J) < 2) or (M(I,J) > 3));
																			boolb := ((cell = '0') and (M(I,J) = 2));
																				boolc := ((cell = '1') and (M(I,J) = 2));
																					boold := (M(I,J) = 3);																			
																						if boold then n := '1'; end if;
																							if boolc then n := '1'; end if;
																								if boola then n := '0'; end if;
																									if boolb then n := '0'; end if;
																										B(I,J) := n;
																											

					
					 
					
						
				
				end loop;
			end loop;
																											decide := 1;
		end if;
																													if decide = 1 and rising_edge(clka) then 
																														for I in 0 to 23 loop
																															for J in 0 to 31 loop
																																A(I,J) := B(I,J);
																															end loop;
																														end loop;
																																	decide := 0;
																													end if;
				
			
			
		
																																		if vidon = '1' then
																																			row := to_integer(unsigned(vcs-vbp));
																																			row := row/20;
																																			col := to_integer(unsigned(hcs-hbp));
																																			col := col/20;
																																			--B(5)(5) := state(bool_1,bool_2,false,bool_4);
																														--					if M(5,5) = 5 then blue <= '1';else blue <= '0'; end if;
																														--						if M(5,5) = 4 then navy <= '1';else navy <= '0'; end if;
																														--							if M(5,5) = 3 then red <= '1';else red <= '0'; end if;
																														--								if M(5,5) = 0 then green <= '1';else green <= '0'; end if;
																																				red <= A(row,col);
																																					--blue <= B(2,2);
																																			--green <= test;
																																			--report "VALUE" & integer'image(test);
--																																			if M(2,1) = 3 then blue <= '1';
--																																				elsif M(7,8) = 3 then green <= '1';
--																																					elsif M(7,1) = 3 then red <= '1';
--																																						elsif M(2,8) = 3 then navy <= '1';
--																																							else green <= '0';red <= '0';blue <= '0';navy <= '0';
																																			--end if;
																																		end if;	
			
--			red <= '0';
--			green <= '0';
--			blue <= '0';
--			if vidon = '1' then
--			red <= vcs(4);-- & vcs(4) & vcs(4);
--			green <= not vcs(4);-- & vcs(4) & vcs(4));
--			end if;
			
	
	end process;

	
end GoL_a;	
	
